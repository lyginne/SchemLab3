@00000000
08 00 00 0C 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
8C 09 00 78 00 00 00 00 AC 09 00 70 42 00 00 10 
8C 08 02 00 00 00 00 00 21 08 00 01 21 08 00 01 
21 08 00 01 21 08 00 01 08 00 00 0E 21 08 00 01 
@00000200
00 00 00 01 00 00 FF FF 
