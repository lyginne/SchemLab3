@00000000
08 00 00 07 00 00 00 00 00 00 00 00 00 00 00 00 
31 08 00 00 31 08 00 00 42 00 00 10 8C 08 02 00 
8C 09 02 00 21 08 00 0B 01 09 40 22 35 08 00 10 
01 09 40 26 01 09 40 2A 01 09 40 20 11 09 FF F7 
00 00 00 00 
@00000200
00 00 00 01 00 00 FF FF 
